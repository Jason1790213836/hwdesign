logic signed 